module ddr2pe_config#(
    )(
    input   clk,
    input   rst,
    
    input           start,
    output  [1 : 0] ddr_working,
    input   [3 : 0] trans_type,
    input   [1 : 0] 
    );
    
endmodule